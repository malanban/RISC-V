module datapath(
	input clk,
	input reset
);
//`include "programm_counter.sv"
//`include "instruction_memory.sv"
//`include "register.sv"
//`include "alu.sv"
//`include "control.sv"
//`include "alu_control.sv"
//`include "memory.sv"
//`include "multiplexor.sv"
//`include "imm_gen.sv"
//`include "instruction.sv"

endmodule 
